module ecc_192bit
    
endmodule